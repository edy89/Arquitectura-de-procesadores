library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

entity im is
    Port ( address : in  STD_LOGIC_VECTOR(31 downto 0);
           rst : in  STD_LOGIC;
           instruction : out  STD_LOGIC_VECTOR(31 downto 0));
end im;

architecture Behavioral of im is
type rom_type is array (63 downto 0) of std_logic_vector (31 downto 0);                 
    signal ROM : rom_type:= ("00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000",
									  "00000000000000000000000000000000","00000000000000000000000000000000"
									  );
									  

    signal rdata : std_logic_vector(31 downto 0);
begin

    --rdata <= ROM(address);

    process (address)
    begin
        if (rst='1') then
				rdata <= ROM(conv_integer("00000000000000000000000000000000"));
        else
				rdata <= ROM(conv_integer(address));
        end if;
    end process;
end Behavioral;