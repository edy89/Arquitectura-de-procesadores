library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity InstructionMemory is
    Port ( rst : in  STD_LOGIC;
           address : in  STD_LOGIC_VECTOR (31 downto 0);
           imout : out  STD_LOGIC_VECTOR (31 downto 0):=(others=>'0'));
end InstructionMemory;
architecture Behavioral of InstructionMemory is
type rom_type is array (63 downto 0) of STD_LOGIC_VECTOR (31 downto 0);                 
	 signal ROM : rom_type:= (
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","00000001000000000000000000000000",
									  "00000001000000000000000000000000","10010000001001001010000000101011",
									  "10100100000001000000000000010001","10100010000100000011111111111010",
									  "10100000000100000010000000000100","00000001000000000000000000000000");
	signal rdata : std_logic_vector (31 downto 0);
begin
	rdata <= ROM(conv_integer(address));
	process (rst,address)
	begin
		  if (rst = '1') then
				imout <= ROM(conv_integer("00000000000000000000000000000000"));
		  else
				imout <= rdata;
		  end if;
	end process;
end Behavioral;