library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity InstructionMemory is
    Port ( rst : in  STD_LOGIC;
           address : in  STD_LOGIC_VECTOR (31 downto 0);
           imout : out  STD_LOGIC_VECTOR (31 downto 0):=(others=>'0'));
end InstructionMemory;
architecture Behavioral of InstructionMemory is
type rom_type is array (63 downto 0) of STD_LOGIC_VECTOR (31 downto 0);                 
	 signal ROM : rom_type:= (
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									 --- "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "00000001000000000000000000000000",
									  "10010000000100000000000000010000",
									  "10000100010000000000000000000001",
									  "10000000101000000010000000000100",
									  "10000001111000000010000000000000",
									  "10100000000000000110000000000011",
									  "10000001111010000010000000000000",
									  "10110011001101000110000000000001",
									  "10110001001010000110000000000010",
									  "10100010000100000010000000000100",
									  "10100000000100000011111111111000",
									  "10000010000100000010000000000101",
									  "00000001000000000000000000000000");
	signal rdata : std_logic_vector (31 downto 0);
begin
	rdata <= ROM(conv_integer(address));
	process (rst,address)
	begin
		  if (rst = '1') then
				imout <= ROM(conv_integer("00000000000000000000000000000000"));
		  else
				imout <= rdata;
		  end if;
	end process;
end Behavioral;